M�nga DVD-filmer anv�nder css.  F�r att se dessa beh�vs ett bibliotek,
libdvdcss.  Debian kan inte distribuera detta p� grund av juridiska
problem, men det finns tillg�ngligt p� andra platser p� internet.  Om
det �r lagligt f�r dig kan du k�ra skriptet
'/usr/share/doc/libdvdread3/examples/install-css.sh' f�r att h�mta och
installera libdvdcss.
